////////////////////////////////////////////////////////////////////////////////
 /*
 FPGA Project Name     : N - Channel Servo Motor Controller
 Top level Entity Name : Servo_Motor_Controller
 Target Device		   : Cyclone V
 
 Code Author           : Shrajan Bhandary
 Date Created          : 08/03/2019 
 Location 			   : University of Leeds
 Module 			   : ELEC5566M FPGA Design for System-on-chip
 
 -------------------------------------------------------------------------------
 
 Description of the Verilog Module: 
	The module is used to control a single SG90 Servo Motor. The servo motor 
	requires an input PWM signal to drive to the required angular position. The 
	PWM signal for the SG90 motor should have a clock period of 20 ms. The 
	desired angular position can be obtained by controlling the ON period (duty
	cycle) of the PWM signal. The duty cycle is can be manually varied by 
	changing the 8 bit inputs connected to 8 different slide switches. The value
	of the duty cycle is latched to the output by using a load signal connected 
	to a push button. The servo motor can be initialised to a default position 
	by pressing the reset push button. The default frequency of the clock is 
	128 kHz.
 
 */
//////////////////////////////////////////////////////////////////////////////// 

module Servo_Motor_Controller # (												// Start of the module.
	
	/* Parameter List of the Servo_Motor_Controller */
	parameter 						DUTY_CYCLE_WIDTH = 8   ,					// The default width is 8-bits ( 0 to 255 ) corresponding to ( -90 to +90 ).
	parameter 						PWM_SIGNAL_WIDTH = 12  ,					// The required width is 12 bits to enclose maximum value of 2560 (20ms) with a clock of 128 kHz frequency.
	parameter						MAX_CLOCK_CYCLES = 2560 					// With a clock of 128 kHz frequency, 2560 clock cycles are required to generate 20 ms.
	
)(	
	/* Port List of the Servo_Motor_Controller */
	input 							CLOCK_SIGNAL      ,							// Connects to the hardware clock to generate the required PWM signal.
	input 							CLOCK_ENABLE      ,							// Servo motor turns only if enable is HIGH.
	input 							SERVO_RESET       ,							// Servo resets to default when reset becomes HIGH.
	input 							LOAD_SIGNAL       ,							// Latch the duty cycle of the PWM signal.
	input  [(DUTY_CYCLE_WIDTH-1):0]	DUTY_CYCLE_CONTROL,							// Controls the duty cycle of the PWM signal, thus controlling the angle.
	output 							PWM_SIGNAL 									// The output of the module that is the input to the Servo motor.
);
	/* Register List of the Servo_Motor_Controller */
	wire [(PWM_SIGNAL_WIDTH-1):0] CURRENT_CLOCK_CYCLES;							// This holds the number of clock cycles generated by the clock with 128 kHz frequency.
	reg  [(PWM_SIGNAL_WIDTH-1):0] REQUIRED_ON_CYCLES  ;							// The ON period (duty cycle) is determined by the 8-bit input.  
	wire DIVIDED_CLOCK_SIGNAL;													// Output of the frequency divider circuit that converts current clock frequency to the default value.
	
	/* Local Parameter List of the Servo_Motor_Controller */
	localparam DEFAULT_ON_CYCLES = {(PWM_SIGNAL_WIDTH){12'd192}}; 				// To set the servo to angle 0, 1.5ms is required which corresponds to 192 clock cycles.
	localparam OFFSET_ON_CYCLES  = {(PWM_SIGNAL_WIDTH){12'd64}} ;				// The on cycles vary from 64(0.5ms) to 320(2.5ms) to turn angles from -90 to 90.
    
	/* Check status of load signal and rest and then take necessary actions */
	always @ ( posedge LOAD_SIGNAL or posedge SERVO_RESET ) 					// Always statement is used to set the required on cycle depending on the value of the 8-bit input.
		begin																	// The sensitivity list contains the latch signal and reset signal.
		
			if ( SERVO_RESET )													// Check if reset is HIGH.
				begin 
					REQUIRED_ON_CYCLES <= DEFAULT_ON_CYCLES;					// Set the servo to its default position if the reset if HIGH.
				end
				
			else if ( CLOCK_ENABLE ) 											// Check if clock enable is HIGH.
				begin
					REQUIRED_ON_CYCLES <= DUTY_CYCLE_CONTROL + OFFSET_ON_CYCLES;// 	Assigning value to the on cycle based upon the duty cycle and the offset.
				end
		end
	
	/* Instantiating N Bit Counter to generate the required clock cycles for the servo motor. */
	N_Bit_Counter #           (															
		. COUNTER_VALUE_WIDTH ( PWM_SIGNAL_WIDTH     ),							// Setting the parameter values.
		. COUNTER_MAX_VALUE   ( MAX_CLOCK_CYCLES     )
		
	) Cycle_Generator         (
		. COUNTER_CLOCK       ( CLOCK_SIGNAL		 ),							// Setting the connections to their corresponding ports. 
		. COUNTER_RESET       ( SERVO_RESET          ),
		. COUNTER_ENABLE      ( CLOCK_ENABLE         ), 
		. COUNTER_VALUE		  ( CURRENT_CLOCK_CYCLES )
	);
	
	/* Instantiating N Bit Comparator to generate the HIGH cycles of the PWM signal. */
	N_Bit_Comparator #    	 (														
		. NUMBER_WIDTH       ( PWM_SIGNAL_WIDTH      )							// Setting the parameter values.
		
	) On_Period_Generator    (
		. FIRST_NUMBER       ( REQUIRED_ON_CYCLES   ),							// Setting the connections to their corresponding ports. 
		. SECOND_NUMBER      ( CURRENT_CLOCK_CYCLES ),
		. FN_GREATER_THAN_SN ( PWM_SIGNAL           ) 
	);
	
endmodule																		// End of the module.